`timescale 1ns / 1ps  

import core_pkg::*;

module IF_to_ID_Reg (
  input logic clk,
  input logic rst_n

  );

endmodule
